/***********************************************************
 * File: Priority_Resolver.v
 * Developer: 
 * Description: 
 ************************************************************/

module Priority_Resolver();

endmodule