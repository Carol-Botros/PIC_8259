/***********************************************************
 * File: TB_In_Service.v
 * Developer: 
 * Description: 
 ************************************************************/

`include "../HDL/In_Service.v"

module TB_In_Service();

endmodule