/***********************************************************
 * File: TB_Cascade_Buffer_Comparator.v
 * Developer: 
 * Description: 
 ************************************************************/

`include "../HDL/Cascade_Buffer_Comparator.v"

module TB_Cascade_Buffer_Comparator();


endmodule