/***********************************************************
 * File: In_Mask_Reg.v
 * Developer: 
 * Description: 
 ************************************************************/

module In_Mask_Reg();

endmodule