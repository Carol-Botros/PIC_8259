/***********************************************************
 * File: TB_Interrupt_Reguest.v
 * Developer: 
 * Description: 
 ************************************************************/

`include "../HDL/Interrupt_Reguest.v"

module TB_Interrupt_Reguest();





endmodule

