/***********************************************************
 * File: Cascade_Buffer_Comparator.v
 * Developer: 
 * Description: 
 ************************************************************/

module Cascade_Buffer_Comparator();




endmodule