/***********************************************************
 * File: Read_Write_Logic.v
 * Developer: 
 * Description: 
 ************************************************************/


module Read_Write_Logic();

endmodule