/***********************************************************
 * File: TB_PIC8259A.v
 * Developer: 
 * Description: 
 ************************************************************/

`include "../HDL/PIC8259A.v"

module TB_PIC8259A();

endmodule