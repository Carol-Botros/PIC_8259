/***********************************************************
 * File: In_Service.v
 * Developer: 
 * Description: 
 ************************************************************/

module In_Service();

endmodule