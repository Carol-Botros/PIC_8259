/***********************************************************
 * File: TB_In_Mask_Reg.v
 * Developer: 
 * Description: 
 ************************************************************/

`include "../HDL/In_Mask_Reg.v"

module TB_In_Mask_Reg();

endmodule