/***********************************************************
 * File: TB_Data_Bus_Buffer.v
 * Developer: 
 * Description: 
 ************************************************************/

`include "../HDL/Data_Bus_Buffer.v"

module TB_Data_Bus_Buffer();

endmodule