/***********************************************************
 * File: Interrupt_Reguest.v
 * Developer: 
 * Description: 
 ************************************************************/

module Interrupt_Reguest();





endmodule

