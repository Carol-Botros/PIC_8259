/***********************************************************
 * File: TB_Read_Write_Logic.v
 * Developer: 
 * Description: 
 ************************************************************/

`include "../HDL/Read_Write_Logic.v"

module TB_Read_Write_Logic();

endmodule