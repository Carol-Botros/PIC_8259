/***********************************************************
 * File: Control_Logic.v
 * Developer: 
 * Description: 
 ************************************************************/

module Control_Logic();

endmodule