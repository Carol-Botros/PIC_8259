/***********************************************************
 * File: TB_Control_Logic.v
 * Developer: 
 * Description: 
 ************************************************************/

`include "../HDL/Control_Logic.v"

module TB_Control_Logic();



endmodule