/***********************************************************
 * File: TB_Priority_Resolver.v
 * Developer: 
 * Description: 
 ************************************************************/

`include "../HDL/Priority_Resolver.v"

module TB_Priority_Resolver();

endmodule