/***********************************************************
 * File: Data_Bus_Buffer.v
 * Developer: 
 * Description: 
 ************************************************************/

module Data_Bus_Buffer();

endmodule