/***********************************************************
 * File: PIC8259A.v
 * Developer: 
 * Description: 
 ************************************************************/

module PIC8259A();

endmodule